o:	Game:@livesi
:
@wordI"corrugated:ET:@letters_foundo:Set:
@hash}I"a;TTF