o:	Game:@livesi:
@wordI"quisling:ET:@letters_foundo:Set:
@hash} F